/*******************************************************************************

-- File Type:    Verilog HDL 
-- Tool Version: VHDL2verilog 20.51
-- Input file was: ..\commonPak.vhd
-- Command line was: D:\SynaptiCAD\bin\win32\vhdl2verilog.exe ..\commonPak.vhd -ncc
-- Date Created: Thu Apr 27 19:58:21 2023

*******************************************************************************/

`define false 1'b 0
`define FALSE 1'b 0
`define true 1'b 1
`define TRUE 1'b 1

