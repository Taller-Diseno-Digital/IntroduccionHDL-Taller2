module tb_contador_regresivo_parametrizable();
logic clk;
logic reset;  
logic a; 
logic y;

