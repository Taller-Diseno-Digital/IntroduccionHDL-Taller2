module topModule(


);


	
ram3 ram_inst(address,clk,data,1'b0,q);