module aletorio();

endmodule